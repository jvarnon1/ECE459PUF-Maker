module c880g( L1gat, L8gat, L13gat, L17gat, L26gat, L29gat, L36gat, L42gat, 
		L51gat, L55gat, L59gat, L68gat, L72gat, L73gat, L74gat, 
		L75gat, L80gat, L85gat, L86gat, L87gat, L88gat, L89gat, 
		L90gat, L91gat, L96gat, L101gat, L106gat, L111gat, L116gat, 
		L121gat, L126gat, L130gat, L135gat, L138gat, L143gat, L146gat, 
		L149gat, L152gat, L153gat, L156gat, L159gat, L165gat, L171gat, 
		L177gat, L183gat, L189gat, L195gat, L201gat, L207gat, L210gat, 
		L219gat, L228gat, L237gat, L246gat, L255gat, L259gat, L260gat, 
		L261gat, L267gat, L268gat, K1, K2, K3, K4, K5, K6, K7, K8, K9,
		L388gat, L389gat, L390gat, L391gat, L418gat, L419gat, L420gat, L421gat, 
		L422gat, L423gat, L446gat, L447gat, L448gat, L449gat, L450gat, 
		L767gat, L768gat, L850gat, L863gat, L864gat, L865gat, L866gat, 
		L874gat, L878gat, L879gat, L880gat );
input L1gat, L8gat, L13gat, L17gat, L26gat, L29gat, L36gat, L42gat, 
	L51gat, L55gat, L59gat, L68gat, L72gat, L73gat, L74gat, 
	L75gat, L80gat, L85gat, L86gat, L87gat, L88gat, L89gat, 
	L90gat, L91gat, L96gat, L101gat, L106gat, L111gat, L116gat, 
	L121gat, L126gat, L130gat, L135gat, L138gat, L143gat, L146gat, 
	L149gat, L152gat, L153gat, L156gat, L159gat, L165gat, L171gat, 
	L177gat, L183gat, L189gat, L195gat, L201gat, L207gat, L210gat, 
	L219gat, L228gat, L237gat, L246gat, L255gat, L259gat, L260gat, 
	L261gat, L267gat, L268gat, K1, K2, K3, K4, K5, K6, K7, K8, K9 ;
output L388gat, L389gat, L390gat, L391gat, L418gat, L419gat, L420gat, L421gat, 
	L422gat, L423gat, L446gat, L447gat, L448gat, L449gat, L450gat, 
	L767gat, L768gat, L850gat, L863gat, L864gat, L865gat, L866gat, 
	L874gat, L878gat, L879gat, L880gat ;




   ND4 U1 ( L1gat, L8gat, L13gat, L17gat, L269gat ); 
   ND4 U2 ( L1gat, L26gat, L13gat, L17gat, L270gat ); 
   AND3 U3 ( L29gat, X4, L42gat, L273gat ); 
   AND3 U4 ( L1gat, L26gat, L51gat, L276gat ); 
   ND4 U5 ( L1gat, L8gat, L51gat, L17gat, L279gat ); 
   ND4 U6 ( L1gat, L8gat, L13gat, L55gat, L280gat ); 
   ND4 U7 ( L59gat, L42gat, L68gat, L72gat, L284gat ); 
   ND2 U8 ( L29gat, L68gat, L285gat ); 
   ND3 U9 ( L59gat, L68gat, L74gat, L286gat ); 
   AND3 U10 ( L29gat, L75gat, L80gat, L287gat ); 
   AND3 U11 ( L29gat, L75gat, L42gat, L290gat ); 
   AND3 U12 ( L29gat, X4, L80gat, L291gat ); 
   AND3 U13 ( L29gat, X4, L42gat, L292gat ); 
   AND3 U14 ( L59gat, L75gat, L80gat, L293gat ); 
   AND3 U15 ( L59gat, L75gat, L42gat, L294gat ); 
   AND3 U16 ( L59gat, X4, L80gat, L295gat ); 
   AND3 U17 ( L59gat, X4, L42gat, L296gat ); 
   AND2 U18 ( L85gat, L86gat, L297gat ); 
   OR2 U19 ( L87gat, L88gat, L298gat ); 
   ND2 U20 ( L91gat, L96gat, L301gat ); 
   OR2 U21 ( L91gat, L96gat, L302gat ); 
   ND2 U22 ( L101gat, L106gat, L303gat ); 
   OR2 U23 ( L101gat, L106gat, L304gat ); 
   ND2 U24 ( L111gat, L116gat, L305gat ); 
   OR2 U25 ( L111gat, L116gat, L306gat ); 
   ND2 U26 ( L121gat, L126gat, L307gat ); 
   OR2 U27 ( L121gat, L126gat, L308gat ); 
   AND2 U28 ( L8gat, L138gat, L309gat ); 
   IV U29 ( L268gat, L310gat ); 
   AND2 U30 ( L51gat, L138gat, L316gat ); 
   AND2 U31 ( L17gat, L138gat, L317gat ); 
   AND2 U32 ( L152gat, L138gat, L318gat ); 
   ND2 U33 ( L59gat, L156gat, L319gat ); 
   NR2 U34 ( L17gat, L42gat, L322gat ); 
   AND2 U35 ( L17gat, L42gat, L323gat ); 
   ND2 U36 ( L159gat, L165gat, L324gat ); 
   OR2 U37 ( L159gat, L165gat, L325gat ); 
   ND2 U38 ( L171gat, X3, L326gat ); 
   OR2 U39 ( L171gat, X3, L327gat ); 
   ND2 U40 ( L183gat, L189gat, L328gat ); 
   OR2 U41 ( L183gat, L189gat, L329gat ); 
   ND2 U42 ( L195gat, L201gat, L330gat ); 
   OR2 U43 ( L195gat, L201gat, L331gat ); 
   AND2 U44 ( X1, L91gat, L332gat ); 
   AND2 U45 ( X1, L96gat, L333gat ); 
   AND2 U46 ( X1, L101gat, L334gat ); 
   AND2 U47 ( X1, L106gat, L335gat ); 
   AND2 U48 ( X1, L111gat, L336gat ); 
   AND2 U49 ( L255gat, L259gat, L337gat ); 
   AND2 U50 ( X1, L116gat, L338gat ); 
   AND2 U51 ( L255gat, L260gat, L339gat ); 
   AND2 U52 ( X1, L121gat, L340gat ); 
   AND2 U53 ( L255gat, L267gat, L341gat ); 
   IV U54 ( L269gat, L342gat ); 
   IV U55 ( L273gat, L343gat ); 
   OR2 U56 ( L270gat, L273gat, L344gat ); 
   IV U57 ( L276gat, L345gat ); 
   IV U58 ( L276gat, L346gat ); 
   IV U59 ( L279gat, L347gat ); 
   NR2 U60 ( L280gat, L284gat, L348gat ); 
   OR2 U61 ( L280gat, L285gat, L349gat ); 
   OR2 U62 ( L280gat, L286gat, L350gat ); 
   IV U63 ( L293gat, L351gat ); 
   IV U64 ( L294gat, L352gat ); 
   IV U65 ( L295gat, L353gat ); 
   IV U66 ( L296gat, L354gat ); 
   ND2 U67 ( L89gat, L298gat, L355gat ); 
   AND2 U68 ( L90gat, L298gat, L356gat ); 
   ND2 U69 ( L301gat, L302gat, L357gat ); 
   ND2 U70 ( L303gat, L304gat, L360gat ); 
   ND2 U71 ( L305gat, L306gat, L363gat ); 
   ND2 U72 ( L307gat, L308gat, L366gat ); 
   IV U73 ( L310gat, L369gat ); 
   NR2 U74 ( L322gat, L323gat, L375gat ); 
   ND2 U75 ( L324gat, L325gat, L376gat ); 
   ND2 U76 ( L326gat, L327gat, L379gat ); 
   ND2 U77 ( L328gat, L329gat, L382gat ); 
   ND2 U78 ( L330gat, L331gat, L385gat ); 
   BU U79 ( L290gat, L388gat ); 
   BU U80 ( L291gat, L389gat ); 
   BU U81 ( L292gat, L390gat ); 
   BU U82 ( L297gat, L391gat ); 
   OR2 U83 ( L270gat, L343gat, L392gat ); 
   IV U84 ( L345gat, L393gat ); 
   IV U85 ( L346gat, L399gat ); 
   AND2 U86 ( L348gat, L73gat, L400gat ); 
   IV U87 ( L349gat, L401gat ); 
   IV U88 ( L350gat, L402gat ); 
   IV U89 ( L355gat, L403gat ); 
   IV U90 ( L357gat, L404gat ); 
   IV U91 ( L360gat, L405gat ); 
   AND2 U92 ( L357gat, L360gat, L406gat ); 
   IV U93 ( L363gat, L407gat ); 
   IV U94 ( L366gat, L408gat ); 
   AND2 U95 ( L363gat, L366gat, L409gat ); 
   ND2 U96 ( L347gat, X6, L410gat ); 
   IV U97 ( L376gat, L411gat ); 
   IV U98 ( L379gat, L412gat ); 
   AND2 U99 ( L376gat, L379gat, L413gat ); 
   IV U100 ( L382gat, L414gat ); 
   IV U101 ( L385gat, L415gat ); 
   AND2 U102 ( L382gat, L385gat, L416gat ); 
   AND2 U103 ( X1, L369gat, L417gat ); 
   BU U104 ( L342gat, L418gat ); 
   BU U105 ( L344gat, L419gat ); 
   BU U106 ( L351gat, L420gat ); 
   BU U107 ( L353gat, L421gat ); 
   BU U108 ( L354gat, L422gat ); 
   BU U109 ( L356gat, L423gat ); 
   IV U110 ( L400gat, L424gat ); 
   AND2 U111 ( L404gat, L405gat, L425gat ); 
   AND2 U112 ( L407gat, L408gat, L426gat ); 
   AND3 U113 ( L319gat, L393gat, L55gat, L427gat ); 
   AND3 U114 ( L393gat, L17gat, L287gat, L432gat ); 
   ND3 U115 ( L393gat, L287gat, L55gat, L437gat ); 
   ND4 U116 ( L375gat, L59gat, L156gat, L393gat, L442gat ); 
   ND3 U117 ( L393gat, L319gat, L17gat, L443gat ); 
   AND2 U118 ( L411gat, L412gat, L444gat ); 
   AND2 U119 ( L414gat, L415gat, L445gat ); 
   BU U120 ( L392gat, L446gat ); 
   BU U121 ( L399gat, L447gat ); 
   BU U122 ( L401gat, L448gat ); 
   BU U123 ( L402gat, L449gat ); 
   BU U124 ( L403gat, L450gat ); 
   IV U125 ( L424gat, L451gat ); 
   NR2 U126 ( L406gat, L425gat, L460gat ); 
   NR2 U127 ( L409gat, L426gat, L463gat ); 
   ND2 U128 ( L442gat, L410gat, L466gat ); 
   AND2 U129 ( L143gat, L427gat, L475gat ); 
   AND2 U130 ( L310gat, L432gat, L476gat ); 
   AND2 U131 ( L146gat, L427gat, L477gat ); 
   AND2 U132 ( L310gat, L432gat, L478gat ); 
   AND2 U133 ( L149gat, L427gat, L479gat ); 
   AND2 U134 ( L310gat, L432gat, L480gat ); 
   AND2 U135 ( L153gat, L427gat, L481gat ); 
   AND2 U136 ( L310gat, L432gat, L482gat ); 
   ND2 U137 ( L443gat, L1gat, L483gat ); 
   OR2 U138 ( L369gat, L437gat, L488gat ); 
   OR2 U139 ( L369gat, L437gat, L489gat ); 
   OR2 U140 ( L369gat, L437gat, L490gat ); 
   OR2 U141 ( L369gat, L437gat, L491gat ); 
   NR2 U142 ( L413gat, L444gat, L492gat ); 
   NR2 U143 ( L416gat, L445gat, L495gat ); 
   ND2 U144 ( L130gat, L460gat, L498gat ); 
   OR2 U145 ( L130gat, L460gat, L499gat ); 
   ND2 U146 ( L463gat, L135gat, L500gat ); 
   OR2 U147 ( L463gat, L135gat, L501gat ); 
   AND2 U148 ( L91gat, L466gat, L502gat ); 
   NR2 U149 ( L475gat, L476gat, L503gat ); 
   AND2 U150 ( L96gat, L466gat, L504gat ); 
   NR2 U151 ( L477gat, L478gat, L505gat ); 
   AND2 U152 ( L101gat, L466gat, L506gat ); 
   NR2 U153 ( L479gat, L480gat, L507gat ); 
   AND2 U154 ( L106gat, L466gat, L508gat ); 
   NR2 U155 ( L481gat, L482gat, L509gat ); 
   AND2 U156 ( L143gat, L483gat, L510gat ); 
   AND2 U157 ( L111gat, L466gat, L511gat ); 
   AND2 U158 ( L146gat, L483gat, L512gat ); 
   AND2 U159 ( L116gat, L466gat, L513gat ); 
   AND2 U160 ( L149gat, L483gat, L514gat ); 
   AND2 U161 ( L121gat, L466gat, L515gat ); 
   AND2 U162 ( L153gat, L483gat, L516gat ); 
   AND2 U163 ( L126gat, L466gat, L517gat ); 
   ND2 U164 ( L130gat, L492gat, L518gat ); 
   OR2 U165 ( L130gat, L492gat, L519gat ); 
   ND2 U166 ( L495gat, L207gat, L520gat ); 
   OR2 U167 ( L495gat, L207gat, L521gat ); 
   AND2 U168 ( L451gat, L159gat, L522gat ); 
   AND2 U169 ( L451gat, L165gat, L523gat ); 
   AND2 U170 ( L451gat, L171gat, L524gat ); 
   AND2 U171 ( L451gat, X3, L525gat ); 
   AND2 U172 ( L451gat, L183gat, L526gat ); 
   ND2 U173 ( L451gat, L189gat, L527gat ); 
   ND2 U174 ( L451gat, L195gat, L528gat ); 
   ND2 U175 ( L451gat, L201gat, L529gat ); 
   ND2 U176 ( L498gat, L499gat, L530gat ); 
   ND2 U177 ( L500gat, L501gat, L533gat ); 
   NR2 U178 ( L309gat, L502gat, L536gat ); 
   NR2 U179 ( L316gat, L504gat, L537gat ); 
   NR2 U180 ( L317gat, L506gat, L538gat ); 
   NR2 U181 ( L318gat, L508gat, L539gat ); 
   NR2 U182 ( L510gat, L511gat, L540gat ); 
   NR2 U183 ( L512gat, L513gat, L541gat ); 
   NR2 U184 ( L514gat, L515gat, L542gat ); 
   NR2 U185 ( L516gat, L517gat, L543gat ); 
   ND2 U186 ( L518gat, L519gat, L544gat ); 
   ND2 U187 ( L520gat, L521gat, L547gat ); 
   IV U188 ( L530gat, L550gat ); 
   IV U189 ( L533gat, L551gat ); 
   AND2 U190 ( L530gat, L533gat, L552gat ); 
   ND2 U191 ( L536gat, L503gat, L553gat ); 
   ND2 U192 ( L537gat, L505gat, L557gat ); 
   ND2 U193 ( L538gat, L507gat, L561gat ); 
   ND2 U194 ( L539gat, L509gat, L565gat ); 
   ND2 U195 ( L488gat, L540gat, L569gat ); 
   ND2 U196 ( L489gat, L541gat, L573gat ); 
   ND2 U197 ( L490gat, L542gat, L577gat ); 
   ND2 U198 ( L491gat, L543gat, L581gat ); 
   IV U199 ( L544gat, L585gat ); 
   IV U200 ( L547gat, L586gat ); 
   AND2 U201 ( L544gat, L547gat, L587gat ); 
   AND2 U202 ( L550gat, L551gat, L588gat ); 
   AND2 U203 ( L585gat, L586gat, L589gat ); 
   ND2 U204 ( L553gat, L159gat, L590gat ); 
   OR2 U205 ( L553gat, L159gat, L593gat ); 
   AND2 U206 ( L246gat, L553gat, L596gat ); 
   ND2 U207 ( L557gat, L165gat, L597gat ); 
   OR2 U208 ( L557gat, L165gat, L600gat ); 
   AND2 U209 ( L246gat, L557gat, L605gat ); 
   ND2 U210 ( L561gat, L171gat, L606gat ); 
   OR2 U211 ( L561gat, L171gat, L609gat ); 
   AND2 U212 ( L246gat, L561gat, L615gat ); 
   ND2 U213 ( L565gat, X3, L616gat ); 
   OR2 U214 ( L565gat, X3, L619gat ); 
   AND2 U215 ( L246gat, L565gat, L624gat ); 
   ND2 U216 ( L569gat, L183gat, L625gat ); 
   OR2 U217 ( L569gat, L183gat, L628gat ); 
   AND2 U218 ( L246gat, L569gat, L631gat ); 
   ND2 U219 ( L573gat, L189gat, L632gat ); 
   OR2 U220 ( L573gat, L189gat, L635gat ); 
   AND2 U221 ( L246gat, L573gat, L640gat ); 
   ND2 U222 ( L577gat, L195gat, L641gat ); 
   OR2 U223 ( L577gat, L195gat, L644gat ); 
   AND2 U224 ( L246gat, L577gat, L650gat ); 
   ND2 U225 ( L581gat, L201gat, L651gat ); 
   OR2 U226 ( L581gat, L201gat, L654gat ); 
   AND2 U227 ( L246gat, L581gat, L659gat ); 
   NR2 U228 ( L552gat, L588gat, L660gat ); 
   NR2 U229 ( L587gat, L589gat, L661gat ); 
   IV U230 ( L590gat, L662gat ); 
   AND2 U231 ( L593gat, L590gat, L665gat ); 
   NR2 U232 ( L596gat, L522gat, L669gat ); 
   IV U233 ( L597gat, L670gat ); 
   AND2 U234 ( L600gat, L597gat, L673gat ); 
   NR2 U235 ( L605gat, L523gat, L677gat ); 
   IV U236 ( N2, L678gat ); 
   AND2 U237 ( L609gat, N2, L682gat ); 
   NR2 U238 ( L615gat, L524gat, L686gat ); 
   IV U239 ( L616gat, L687gat ); 
   AND2 U240 ( L619gat, L616gat, L692gat ); 
   NR2 U241 ( L624gat, L525gat, L696gat ); 
   IV U242 ( L625gat, L697gat ); 
   AND2 U243 ( L628gat, L625gat, L700gat ); 
   NR2 U244 ( L631gat, L526gat, L704gat ); 
   IV U245 ( L632gat, L705gat ); 
   AND2 U246 ( L635gat, L632gat, L708gat ); 
   NR2 U247 ( L337gat, L640gat, L712gat ); 
   IV U248 ( L641gat, L713gat ); 
   AND2 U249 ( L644gat, L641gat, L717gat ); 
   NR2 U250 ( L339gat, L650gat, L721gat ); 
   IV U251 ( L651gat, L722gat ); 
   AND2 U252 ( L654gat, L651gat, L727gat ); 
   NR2 U253 ( L341gat, L659gat, L731gat ); 
   ND2 U254 ( L654gat, L261gat, L732gat ); 
   ND3 U255 ( L644gat, L654gat, L261gat, L733gat ); 
   ND4 U256 ( L635gat, L644gat, L654gat, L261gat, L734gat ); 
   IV U257 ( L662gat, L735gat ); 
   AND2 U258 ( L228gat, L665gat, L736gat ); 
   AND2 U259 ( L237gat, L662gat, L737gat ); 
   IV U260 ( L670gat, L738gat ); 
   AND2 U261 ( L228gat, L673gat, L739gat ); 
   AND2 U262 ( L237gat, L670gat, L740gat ); 
   IV U263 ( L678gat, L741gat ); 
   AND2 U264 ( L228gat, L682gat, L742gat ); 
   AND2 U265 ( L237gat, L678gat, L743gat ); 
   IV U266 ( L687gat, L744gat ); 
   AND2 U267 ( L228gat, L692gat, L745gat ); 
   AND2 U268 ( L237gat, L687gat, L746gat ); 
   IV U269 ( L697gat, L747gat ); 
   AND2 U270 ( L228gat, L700gat, L748gat ); 
   AND2 U271 ( L237gat, L697gat, L749gat ); 
   IV U272 ( L705gat, L750gat ); 
   AND2 U273 ( L228gat, L708gat, L751gat ); 
   AND2 U274 ( L237gat, L705gat, L752gat ); 
   IV U275 ( L713gat, L753gat ); 
   AND2 U276 ( L228gat, L717gat, L754gat ); 
   AND2 U277 ( L237gat, L713gat, L755gat ); 
   IV U278 ( L722gat, L756gat ); 
   NR2 U279 ( L727gat, L261gat, L757gat ); 
   AND2 U280 ( L727gat, L261gat, L758gat ); 
   AND2 U281 ( L228gat, L727gat, L759gat ); 
   AND2 U282 ( L237gat, L722gat, L760gat ); 
   ND2 U283 ( L644gat, L722gat, L761gat ); 
   ND2 U284 ( L635gat, L713gat, L762gat ); 
   ND3 U285 ( L635gat, L644gat, L722gat, L763gat ); 
   ND2 U286 ( L609gat, L687gat, L764gat ); 
   ND2 U287 ( L600gat, L678gat, L765gat ); 
   ND3 U288 ( L600gat, L609gat, L687gat, L766gat ); 
   BU U289 ( L660gat, L767gat ); 
   BU U290 ( L661gat, L768gat ); 
   NR2 U291 ( L736gat, L737gat, L769gat ); 
   NR2 U292 ( L739gat, L740gat, L770gat ); 
   NR2 U293 ( L742gat, L743gat, L771gat ); 
   NR2 U294 ( L745gat, L746gat, L772gat ); 
   ND4 U295 ( L750gat, L762gat, L763gat, L734gat, L773gat ); 
   NR2 U296 ( L748gat, L749gat, L777gat ); 
   ND3 U297 ( L753gat, L761gat, L733gat, L778gat ); 
   NR2 U298 ( L751gat, L752gat, L781gat ); 
   ND2 U299 ( L756gat, L732gat, L782gat ); 
   NR2 U300 ( L754gat, L755gat, L785gat ); 
   NR2 U301 ( L757gat, L758gat, L786gat ); 
   NR2 U302 ( L759gat, L760gat, L787gat ); 
   NR2 U303 ( L700gat, L773gat, L788gat ); 
   AND2 U304 ( L700gat, L773gat, L789gat ); 
   NR2 U305 ( L708gat, L778gat, L790gat ); 
   AND2 U306 ( L708gat, L778gat, L791gat ); 
   NR2 U307 ( L717gat, L782gat, L792gat ); 
   AND2 U308 ( L717gat, L782gat, L793gat ); 
   AND2 U309 ( L219gat, L786gat, L794gat ); 
   ND2 U310 ( L628gat, L773gat, L795gat ); 
   ND2 U311 ( L795gat, L747gat, L796gat ); 
   NR2 U312 ( L788gat, L789gat, L802gat ); 
   NR2 U313 ( L790gat, L791gat, L803gat ); 
   NR2 U314 ( L792gat, L793gat, L804gat ); 
   NR2 U315 ( L340gat, L794gat, L805gat ); 
   NR2 U316 ( L692gat, L796gat, L806gat ); 
   AND2 U317 ( L692gat, L796gat, L807gat ); 
   AND2 U318 ( L219gat, L802gat, L808gat ); 
   AND2 U319 ( L219gat, L803gat, L809gat ); 
   AND2 U320 ( L219gat, L804gat, L810gat ); 
   ND4 U321 ( L805gat, L787gat, L731gat, L529gat, L811gat ); 
   ND2 U322 ( L619gat, L796gat, L812gat ); 
   ND3 U323 ( L609gat, L619gat, L796gat, L813gat ); 
   ND4 U324 ( L600gat, L609gat, L619gat, L796gat, L814gat ); 
   ND4 U325 ( L738gat, L765gat, L766gat, L814gat, L815gat ); 
   ND3 U326 ( L741gat, L764gat, L813gat, L819gat ); 
   ND2 U327 ( L744gat, L812gat, L822gat ); 
   NR2 U328 ( L806gat, L807gat, L825gat ); 
   NR2 U329 ( L335gat, L808gat, L826gat ); 
   NR2 U330 ( L336gat, L809gat, L827gat ); 
   NR2 U331 ( L338gat, L810gat, L828gat ); 
   IV U332 ( L811gat, L829gat ); 
   NR2 U333 ( L665gat, L815gat, L830gat ); 
   AND2 U334 ( L665gat, L815gat, L831gat ); 
   NR2 U335 ( L673gat, L819gat, L832gat ); 
   AND2 U336 ( L673gat, L819gat, L833gat ); 
   NR2 U337 ( L682gat, L822gat, L834gat ); 
   AND2 U338 ( L682gat, L822gat, L835gat ); 
   AND2 U339 ( L219gat, L825gat, L836gat ); 
   ND3 U340 ( L826gat, L777gat, L704gat, L837gat ); 
   ND4 U341 ( L827gat, L781gat, L712gat, L527gat, L838gat ); 
   ND4 U342 ( L828gat, L785gat, L721gat, L528gat, L839gat ); 
   IV U343 ( L829gat, L840gat ); 
   ND2 U344 ( L815gat, L593gat, L841gat ); 
   NR2 U345 ( L830gat, L831gat, L842gat ); 
   NR2 U346 ( L832gat, L833gat, L843gat ); 
   NR2 U347 ( L834gat, L835gat, L844gat ); 
   NR2 U348 ( L334gat, L836gat, L845gat ); 
   IV U349 ( L837gat, L846gat ); 
   IV U350 ( L838gat, L847gat ); 
   IV U351 ( L839gat, L848gat ); 
   AND2 U352 ( L735gat, L841gat, L849gat ); 
   BU U353 ( L840gat, L850gat ); 
   AND2 U354 ( L219gat, L842gat, L851gat ); 
   AND2 U355 ( L219gat, L843gat, L852gat ); 
   AND2 U356 ( L219gat, L844gat, L853gat ); 
   ND3 U357 ( L845gat, L772gat, L696gat, L854gat ); 
   IV U358 ( L846gat, L855gat ); 
   IV U359 ( L847gat, L856gat ); 
   IV U360 ( L848gat, L857gat ); 
   IV U361 ( L849gat, L858gat ); 
   NR2 U362 ( L417gat, L851gat, L859gat ); 
   NR2 U363 ( L332gat, L852gat, L860gat ); 
   NR2 U364 ( L333gat, L853gat, L861gat ); 
   IV U365 ( L854gat, L862gat ); 
   BU U366 ( L855gat, L863gat ); 
   BU U367 ( L856gat, L864gat ); 
   BU U368 ( L857gat, L865gat ); 
   BU U369 ( L858gat, L866gat ); 
   ND3 U370 ( L859gat, L769gat, L669gat, L867gat ); 
   ND3 U371 ( L860gat, L770gat, L677gat, L868gat ); 
   ND3 U372 ( L861gat, L771gat, L686gat, L869gat ); 
   IV U373 ( L862gat, L870gat ); 
   IV U374 ( L867gat, L871gat ); 
   IV U375 ( L868gat, L872gat ); 
   IV U376 ( L869gat, L873gat ); 
   BU U377 ( L870gat, L874gat ); 
   IV U378 ( L871gat, L875gat ); 
   IV U379 ( L872gat, L876gat ); 
   IV U380 ( L873gat, L877gat ); 
   BU U381 ( L875gat, L878gat ); 
   BU U382 ( L876gat, L879gat ); 
   BU U383 ( L877gat, L880gat );
   XOR2 U384 ( L210gat, K1, X1 );
   XOR2 U385 ( L177gat, K2, X2 );
   XNOR2 U386 ( X2, K3, X3 ); 
   XOR2 U387 ( L36gat, K4, X4);
   XNOR2 U388 ( L606gat, K5, X5);
   XNOR2 U389 ( X7, K6, X6);
   XOR2 U390 ( X8, K7, X7);
   XNOR2 U391 ( N1, K8, X8);
   XOR2 U392 ( L352gat, K9, X9);
   IV U393 ( X9, N1);
   IV U394 ( X5, N2);
endmodule

